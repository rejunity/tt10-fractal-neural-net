`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a VCD file. You can view it with gtkwave or surfer.
  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, tb);
    #1;
  end

  wire [15:0] out = { {3{uio_out[7]}}, uio_out[6:2], uo_out[7:0] };

`ifndef GL_TEST
  wire [31:0] pop32_data;
  wire [5:0] pop32_count;
  PopCount32 test_pop32(.data(pop32_data), .count(pop32_count));

  wire [63:0] pop64_data;
  wire [6:0] pop64_count;
  PopCount64 test_pop64(.data(pop64_data), .count(pop64_count));

  wire [127:0] pop128_data;
  wire [7:0] pop128_count;
  PopCount128 test_pop128(.data(pop128_data), .count(pop128_count));

`endif

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;
`ifdef GL_TEST
  wire VPWR = 1'b1;
  wire VGND = 1'b0;
`endif

  // Replace tt_um_example with your module name:
  tt_um_rejunity_ternary_dot ternary_dot (

      // Include power ports for the Gate Level test:
`ifdef GL_TEST
      .VPWR(VPWR),
      .VGND(VGND),
`endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

endmodule
